library ieee;
use ieee.std_logic_1164.all;

package LogPackage is

    -- Return ceil(log2(N))
    function log2(N : natural) return natural;

end package LogPackage;

package body LogPackage is

    function log2(N : natural) return natural is
    begin
        if N <= 1 then 
            return 0;
        elsif N <= 2 then 
            return 1;
        elsif N <= 4 then 
            return 2;
        elsif N <= 8 then 
            return 3;
        elsif N <= 16 then 
            return 4;
        elsif N <= 32 then 
            return 5;
        elsif N <= 64 then 
            return 6;
        elsif N <= 128 then 
            return 7;
        else
            return 8;  -- Extend as needed
        end if;
    end function;

end package body LogPackage;
