CONFIGURATION Config_CombMux2_CondS OF ExecUnitTB IS
  FOR Testing
    FOR DUT : TestUnit
      USE ENTITY work.ExecUnit(CombMux2_CondS);
    END FOR;
  END FOR;
END CONFIGURATION Config_CombMux2_CondS;